module decode
//-----------------------------------------------------------------
// Params
//-----------------------------------------------------------------
#(
     parameter SUPPORT_MULDIV   = 1
    ,parameter EXTRA_DECODE_STAGE = 0
)
//-----------------------------------------------------------------
// Ports
//-----------------------------------------------------------------
(
    // Inputs
     input           clk_i
    ,input           rst_i
    ,input           fetch_in_valid_i
    ,input  [127:0]  fetch_in_instr_i
    ,input  [  1:0]  fetch_in_pred_branch_i
    ,input           fetch_in_fault_fetch_i
    ,input           fetch_in_fault_page_i
    ,input  [ 31:0]  fetch_in_pc_i
    ,input           fetch_out0_accept_i
    ,input           fetch_out1_accept_i
    ,input           fetch_out2_accept_i
    ,input           fetch_out3_accept_i
    ,input           branch_request_i
    ,input  [ 31:0]  branch_pc_i
    ,input  [  1:0]  branch_priv_i

    // Outputs
    ,output          fetch_in_accept_o
    ,output          fetch_out0_valid_o
    ,output [ 31:0]  fetch_out0_instr_o
    ,output [ 31:0]  fetch_out0_pc_o
    ,output          fetch_out0_fault_fetch_o
    ,output          fetch_out0_fault_page_o
    ,output          fetch_out0_instr_exec_o
    ,output          fetch_out0_instr_lsu_o
    ,output          fetch_out0_instr_branch_o
    ,output          fetch_out0_instr_mul_o
    ,output          fetch_out0_instr_div_o
    ,output          fetch_out0_instr_csr_o
    ,output          fetch_out0_instr_rd_valid_o
    ,output          fetch_out0_instr_invalid_o
    ,output          fetch_out1_valid_o
    ,output [ 31:0]  fetch_out1_instr_o
    ,output [ 31:0]  fetch_out1_pc_o
    ,output          fetch_out1_fault_fetch_o
    ,output          fetch_out1_fault_page_o
    ,output          fetch_out1_instr_exec_o
    ,output          fetch_out1_instr_lsu_o
    ,output          fetch_out1_instr_branch_o
    ,output          fetch_out1_instr_mul_o
    ,output          fetch_out1_instr_div_o
    ,output          fetch_out1_instr_csr_o
    ,output          fetch_out1_instr_rd_valid_o
    ,output          fetch_out1_instr_invalid_o
    // Outputs for 3rd instruction in fetch bundle (if present)
    ,output          fetch_out2_valid_o
    ,output [ 31:0]  fetch_out2_instr_o
    ,output [ 31:0]  fetch_out2_pc_o
    ,output          fetch_out2_fault_fetch_o
    ,output          fetch_out2_fault_page_o
    ,output          fetch_out2_instr_exec_o
    ,output          fetch_out2_instr_lsu_o
    ,output          fetch_out2_instr_branch_o
    ,output          fetch_out2_instr_mul_o
    ,output          fetch_out2_instr_div_o
    ,output          fetch_out2_instr_csr_o
    ,output          fetch_out2_instr_rd_valid_o
    ,output          fetch_out2_instr_invalid_o
    // Outputs for 4th instruction in fetch bundle (if present)
    ,output          fetch_out3_valid_o
    ,output [ 31:0]  fetch_out3_instr_o
    ,output [ 31:0]  fetch_out3_pc_o
    ,output          fetch_out3_fault_fetch_o
    ,output          fetch_out3_fault_page_o
    ,output          fetch_out3_instr_exec_o
    ,output          fetch_out3_instr_lsu_o
    ,output          fetch_out3_instr_branch_o
    ,output          fetch_out3_instr_mul_o
    ,output          fetch_out3_instr_div_o
    ,output          fetch_out3_instr_csr_o
    ,output          fetch_out3_instr_rd_valid_o
    ,output          fetch_out3_instr_invalid_o
);



wire        enable_muldiv_w     = SUPPORT_MULDIV;

//-----------------------------------------------------------------
// 2 cycle frontend latency
//-----------------------------------------------------------------
generate
if (EXTRA_DECODE_STAGE)
begin
    wire        fetch_in_fault_page_w;
    wire        fetch_in_fault_fetch_w;
    wire [1:0]  fetch_in_pred_branch_w;
    wire [127:0] fetch_in_instr_raw_w;
    wire [127:0] fetch_in_instr_w;
    wire [31:0] fetch_in_pc_w;
    wire        fetch_in_valid_w;

    reg [164:0] fetch_buffer_q;

    always @ (posedge clk_i or posedge rst_i)
    if (rst_i)
        fetch_buffer_q <= 165'b0;
    else if (branch_request_i)
        fetch_buffer_q <= 165'b0;
    else if (!fetch_in_valid_w || fetch_in_accept_o)
        fetch_buffer_q <= {fetch_in_fault_page_i, fetch_in_fault_fetch_i, fetch_in_pred_branch_i, fetch_in_instr_i, fetch_in_pc_i, fetch_in_valid_i};

    assign {fetch_in_fault_page_w, 
            fetch_in_fault_fetch_w, 
            fetch_in_pred_branch_w, 
            fetch_in_instr_raw_w, 
            fetch_in_pc_w, 
            fetch_in_valid_w} = fetch_buffer_q;

    assign fetch_in_instr_w = (fetch_in_fault_page_w | fetch_in_fault_fetch_w) ? 128'b0 : fetch_in_instr_raw_w;

    wire [7:0] info0_in_w;
    wire [9:0] info0_out_w;
    wire [7:0] info1_in_w;
    wire [9:0] info1_out_w;
    wire [7:0] info2_in_w;
    wire [9:0] info2_out_w;
    wire [7:0] info3_in_w;
    wire [9:0] info3_out_w;


    decoder
    u_dec0
    (
         .valid_i(fetch_in_valid_w)
        ,.fetch_fault_i(fetch_in_fault_fetch_w | fetch_in_fault_page_w)
        ,.enable_muldiv_i(enable_muldiv_w)
        ,.opcode_i(fetch_in_instr_w[31:0])

        ,.invalid_o(info0_in_w[7])
        ,.exec_o(info0_in_w[6])
        ,.lsu_o(info0_in_w[5])
        ,.branch_o(info0_in_w[4])
        ,.mul_o(info0_in_w[3])
        ,.div_o(info0_in_w[2])
        ,.csr_o(info0_in_w[1])
        ,.rd_valid_o(info0_in_w[0])
    );

    decoder
    u_dec1
    (
         .valid_i(fetch_in_valid_w)
        ,.fetch_fault_i(fetch_in_fault_fetch_w | fetch_in_fault_page_w)
        ,.enable_muldiv_i(enable_muldiv_w)
        ,.opcode_i(fetch_in_instr_w[63:32])

        ,.invalid_o(info1_in_w[7])
        ,.exec_o(info1_in_w[6])
        ,.lsu_o(info1_in_w[5])
        ,.branch_o(info1_in_w[4])
        ,.mul_o(info1_in_w[3])
        ,.div_o(info1_in_w[2])
        ,.csr_o(info1_in_w[1])
        ,.rd_valid_o(info1_in_w[0])
    );

    decoder
    u_dec2
    (
         .valid_i(fetch_in_valid_w)
        ,.fetch_fault_i(fetch_in_fault_fetch_w | fetch_in_fault_page_w)
        ,.enable_muldiv_i(enable_muldiv_w)
        ,.opcode_i(fetch_in_instr_w[95:64])

        ,.invalid_o(info2_in_w[7])
        ,.exec_o(info2_in_w[6])
        ,.lsu_o(info2_in_w[5])
        ,.branch_o(info2_in_w[4])
        ,.mul_o(info2_in_w[3])
        ,.div_o(info2_in_w[2])
        ,.csr_o(info2_in_w[1])
        ,.rd_valid_o(info2_in_w[0])
    );

    decoder
    u_dec3
    (
         .valid_i(fetch_in_valid_w)
        ,.fetch_fault_i(fetch_in_fault_fetch_w | fetch_in_fault_page_w)
        ,.enable_muldiv_i(enable_muldiv_w)
        ,.opcode_i(fetch_in_instr_w[127:96])

        ,.invalid_o(info3_in_w[7])
        ,.exec_o(info3_in_w[6])
        ,.lsu_o(info3_in_w[5])
        ,.branch_o(info3_in_w[4])
        ,.mul_o(info3_in_w[3])
        ,.div_o(info3_in_w[2])
        ,.csr_o(info3_in_w[1])
        ,.rd_valid_o(info3_in_w[0])
    );

    fetch_fifo
    #( .OPC_INFO_W(10) )
    u_fifo
    (
         .clk_i(clk_i)
        ,.rst_i(rst_i)

        ,.flush_i(branch_request_i)

        // Input side
        ,.push_i(fetch_in_valid_w)
        ,.pc_in_i(fetch_in_pc_w)
        ,.pred_in_i(fetch_in_pred_branch_w)
        ,.data_in_i(fetch_in_instr_w)
        ,.info0_in_i({info0_in_w, fetch_in_fault_page_w, fetch_in_fault_fetch_w})
        ,.info1_in_i({info1_in_w, fetch_in_fault_page_w, fetch_in_fault_fetch_w})
        ,.info2_in_i({info2_in_w, fetch_in_fault_page_w, fetch_in_fault_fetch_w})
        ,.info3_in_i({info3_in_w, fetch_in_fault_page_w, fetch_in_fault_fetch_w})
        ,.accept_o(fetch_in_accept_o)

        // Outputs
        ,.valid0_o(fetch_out0_valid_o)
        ,.pc0_out_o(fetch_out0_pc_o)
        ,.data0_out_o(fetch_out0_instr_o)
        ,.info0_out_o({fetch_out0_instr_invalid_o, fetch_out0_instr_exec_o,
                       fetch_out0_instr_lsu_o,     fetch_out0_instr_branch_o,
                       fetch_out0_instr_mul_o,     fetch_out0_instr_div_o,
                       fetch_out0_instr_csr_o,     fetch_out0_instr_rd_valid_o,
                       fetch_out0_fault_page_o,    fetch_out0_fault_fetch_o})
        ,.pop0_i(fetch_out0_accept_i)

        ,.valid1_o(fetch_out1_valid_o)
        ,.pc1_out_o(fetch_out1_pc_o)
        ,.data1_out_o(fetch_out1_instr_o)
        ,.info1_out_o({fetch_out1_instr_invalid_o, fetch_out1_instr_exec_o,
                       fetch_out1_instr_lsu_o,     fetch_out1_instr_branch_o,
                       fetch_out1_instr_mul_o,     fetch_out1_instr_div_o,
                       fetch_out1_instr_csr_o,     fetch_out1_instr_rd_valid_o,
                       fetch_out1_fault_page_o,    fetch_out1_fault_fetch_o})
        ,.pop1_i(fetch_out1_accept_i)

        ,.valid2_o(fetch_out2_valid_o)
        ,.pc2_out_o(fetch_out2_pc_o)
        ,.data2_out_o(fetch_out2_instr_o)
        ,.info2_out_o({fetch_out2_instr_invalid_o, fetch_out2_instr_exec_o,
                       fetch_out2_instr_lsu_o,     fetch_out2_instr_branch_o,
                       fetch_out2_instr_mul_o,     fetch_out2_instr_div_o,
                       fetch_out2_instr_csr_o,     fetch_out2_instr_rd_valid_o,
                       fetch_out2_fault_page_o,    fetch_out2_fault_fetch_o})
        ,.pop2_i(fetch_out2_accept_i)

        ,.valid3_o(fetch_out3_valid_o)
        ,.pc3_out_o(fetch_out3_pc_o)
        ,.data3_out_o(fetch_out3_instr_o)
        ,.info3_out_o({fetch_out3_instr_invalid_o, fetch_out3_instr_exec_o,
                       fetch_out3_instr_lsu_o,     fetch_out3_instr_branch_o,
                       fetch_out3_instr_mul_o,     fetch_out3_instr_div_o,
                       fetch_out3_instr_csr_o,     fetch_out3_instr_rd_valid_o,
                       fetch_out3_fault_page_o,    fetch_out3_fault_fetch_o})
        ,.pop3_i(fetch_out3_accept_i)
    );
end
//-----------------------------------------------------------------
// 1 cycle frontend latency
//-----------------------------------------------------------------
else
begin
    fetch_fifo
    #( .OPC_INFO_W(2) )
    u_fifo
    (
         .clk_i(clk_i)
        ,.rst_i(rst_i)

        ,.flush_i(branch_request_i)

        // Input side
        ,.push_i(fetch_in_valid_i)
        ,.pc_in_i(fetch_in_pc_i)
        ,.pred_in_i(fetch_in_pred_branch_i)
        ,.data_in_i((fetch_in_fault_page_i | fetch_in_fault_fetch_i) ? 128'b0 : fetch_in_instr_i)
        ,.info0_in_i({fetch_in_fault_page_i, fetch_in_fault_fetch_i})
        ,.info1_in_i({fetch_in_fault_page_i, fetch_in_fault_fetch_i})
        ,.info2_in_i({fetch_in_fault_page_i, fetch_in_fault_fetch_i})
        ,.info3_in_i({fetch_in_fault_page_i, fetch_in_fault_fetch_i})
        ,.accept_o(fetch_in_accept_o)

        // Outputs
        ,.valid0_o(fetch_out0_valid_o)
        ,.pc0_out_o(fetch_out0_pc_o)
        ,.data0_out_o(fetch_out0_instr_o)
        ,.info0_out_o({fetch_out0_fault_page_o, fetch_out0_fault_fetch_o})
        ,.pop0_i(fetch_out0_accept_i)

        ,.valid1_o(fetch_out1_valid_o)
        ,.pc1_out_o(fetch_out1_pc_o)
        ,.data1_out_o(fetch_out1_instr_o)
        ,.info1_out_o({fetch_out1_fault_page_o, fetch_out1_fault_fetch_o})
        ,.pop1_i(fetch_out1_accept_i)

        ,.valid2_o(fetch_out2_valid_o)
        ,.pc2_out_o(fetch_out2_pc_o)
        ,.data2_out_o(fetch_out2_instr_o)
        ,.info2_out_o({fetch_out2_fault_page_o, fetch_out2_fault_fetch_o})
        ,.pop2_i(fetch_out2_accept_i)

        ,.valid3_o(fetch_out3_valid_o)
        ,.pc3_out_o(fetch_out3_pc_o)
        ,.data3_out_o(fetch_out3_instr_o)
        ,.info3_out_o({fetch_out3_fault_page_o, fetch_out3_fault_fetch_o})
        ,.pop3_i(fetch_out3_accept_i)
    );

    decoder
    u_dec0
    (
         .valid_i(fetch_out0_valid_o)
        ,.fetch_fault_i(fetch_out0_fault_fetch_o | fetch_out0_fault_page_o)
        ,.enable_muldiv_i(enable_muldiv_w)
        ,.opcode_i(fetch_out0_instr_o)

        ,.invalid_o(fetch_out0_instr_invalid_o)
        ,.exec_o(fetch_out0_instr_exec_o)
        ,.lsu_o(fetch_out0_instr_lsu_o)
        ,.branch_o(fetch_out0_instr_branch_o)
        ,.mul_o(fetch_out0_instr_mul_o)
        ,.div_o(fetch_out0_instr_div_o)
        ,.csr_o(fetch_out0_instr_csr_o)
        ,.rd_valid_o(fetch_out0_instr_rd_valid_o)
    );

    decoder
    u_dec1
    (
         .valid_i(fetch_out1_valid_o)
        ,.fetch_fault_i(fetch_out1_fault_fetch_o | fetch_out1_fault_page_o)
        ,.enable_muldiv_i(enable_muldiv_w)
        ,.opcode_i(fetch_out1_instr_o)

        ,.invalid_o(fetch_out1_instr_invalid_o)
        ,.exec_o(fetch_out1_instr_exec_o)
        ,.lsu_o(fetch_out1_instr_lsu_o)
        ,.branch_o(fetch_out1_instr_branch_o)
        ,.mul_o(fetch_out1_instr_mul_o)
        ,.div_o(fetch_out1_instr_div_o)
        ,.csr_o(fetch_out1_instr_csr_o)
        ,.rd_valid_o(fetch_out1_instr_rd_valid_o)
    );

    decoder
    u_dec2
    (
         .valid_i(fetch_out2_valid_o)
        ,.fetch_fault_i(fetch_out2_fault_fetch_o | fetch_out2_fault_page_o)
        ,.enable_muldiv_i(enable_muldiv_w)
        ,.opcode_i(fetch_out2_instr_o)

        ,.invalid_o(fetch_out2_instr_invalid_o)
        ,.exec_o(fetch_out2_instr_exec_o)
        ,.lsu_o(fetch_out2_instr_lsu_o)
        ,.branch_o(fetch_out2_instr_branch_o)
        ,.mul_o(fetch_out2_instr_mul_o)
        ,.div_o(fetch_out2_instr_div_o)
        ,.csr_o(fetch_out2_instr_csr_o)
        ,.rd_valid_o(fetch_out2_instr_rd_valid_o)
    );

    decoder
    u_dec3
    (
         .valid_i(fetch_out3_valid_o)
        ,.fetch_fault_i(fetch_out3_fault_fetch_o | fetch_out3_fault_page_o)
        ,.enable_muldiv_i(enable_muldiv_w)
        ,.opcode_i(fetch_out3_instr_o)

        ,.invalid_o(fetch_out3_instr_invalid_o)
        ,.exec_o(fetch_out3_instr_exec_o)
        ,.lsu_o(fetch_out3_instr_lsu_o)
        ,.branch_o(fetch_out3_instr_branch_o)
        ,.mul_o(fetch_out3_instr_mul_o)
        ,.div_o(fetch_out3_instr_div_o)
        ,.csr_o(fetch_out3_instr_csr_o)
        ,.rd_valid_o(fetch_out3_instr_rd_valid_o)
    );
end
endgenerate

endmodule

module fetch_fifo
//-----------------------------------------------------------------
// Params
//-----------------------------------------------------------------
#(
    parameter WIDTH   = 128,
    parameter DEPTH   = 2,
    parameter ADDR_W  = 1,
    parameter OPC_INFO_W = 10
)
//-----------------------------------------------------------------
// Ports
//-----------------------------------------------------------------
(
     input                  clk_i
    ,input                  rst_i

    ,input                  flush_i

    // Input side
    ,input                  push_i
    ,input  [31:0]          pc_in_i
    ,input  [1:0]           pred_in_i
    ,input  [WIDTH-1:0]     data_in_i
    ,input [OPC_INFO_W-1:0] info0_in_i
    ,input [OPC_INFO_W-1:0] info1_in_i
    ,input [OPC_INFO_W-1:0] info2_in_i
    ,input [OPC_INFO_W-1:0] info3_in_i
    ,output                 accept_o

    // Outputs
    ,output                 valid0_o
    ,output  [31:0]         pc0_out_o
    ,output [(WIDTH/4)-1:0] data0_out_o
    ,output[OPC_INFO_W-1:0] info0_out_o
    ,input                  pop0_i

    ,output                 valid1_o
    ,output  [31:0]         pc1_out_o
    ,output [(WIDTH/4)-1:0] data1_out_o
    ,output[OPC_INFO_W-1:0] info1_out_o
    ,input                  pop1_i

    ,output                 valid2_o
    ,output  [31:0]         pc2_out_o
    ,output [(WIDTH/4)-1:0] data2_out_o
    ,output[OPC_INFO_W-1:0] info2_out_o
    ,input                  pop2_i

    ,output                 valid3_o
    ,output  [31:0]         pc3_out_o
    ,output [(WIDTH/4)-1:0] data3_out_o
    ,output[OPC_INFO_W-1:0] info3_out_o
    ,input                  pop3_i
);

//-----------------------------------------------------------------
// Local Params
//-----------------------------------------------------------------
localparam COUNT_W = ADDR_W + 1;

//-----------------------------------------------------------------
// Registers
//-----------------------------------------------------------------
reg [31:0]           pc_q[DEPTH-1:0];
reg                  valid0_q[DEPTH-1:0];
reg                  valid1_q[DEPTH-1:0];
reg                  valid2_q[DEPTH-1:0];
reg                  valid3_q[DEPTH-1:0];
reg [OPC_INFO_W-1:0] info0_q[DEPTH-1:0];
reg [OPC_INFO_W-1:0] info1_q[DEPTH-1:0];
reg [OPC_INFO_W-1:0] info2_q[DEPTH-1:0];
reg [OPC_INFO_W-1:0] info3_q[DEPTH-1:0];
reg [WIDTH-1:0]      ram_q[DEPTH-1:0];
reg [ADDR_W-1:0]     rd_ptr_q;
reg [ADDR_W-1:0]     wr_ptr_q;
reg [COUNT_W-1:0]    count_q;

//-----------------------------------------------------------------
// Sequential
//-----------------------------------------------------------------
wire push_w         = (push_i & accept_o);
wire pop0_w         = (pop0_i & valid0_o);
wire pop1_w         = (pop1_i & valid1_o);
wire pop2_w         = (pop2_i & valid2_o);
wire pop3_w         = (pop3_i & valid3_o);
wire pop_complete_w = (pop0_w | ~valid0_o) & 
                      (pop1_w | ~valid1_o) & 
                      (pop2_w | ~valid2_o) & 
                      (pop3_w | ~valid3_o) &
                      (count_q != 0);
// wire pop_complete_w = ((pop0_w && ~valid1_o) || (pop0_w && ~valid2_o) || (pop0_w && ~valid3_o) || 
//                        (pop1_w && ~valid0_o) || (pop1_w && ~valid2_o) || (pop1_w && ~valid3_o) ||
//                        (pop2_w && ~valid0_o) || (pop2_w && ~valid1_o) || (pop2_w && ~valid3_o) ||
//                        (pop3_w && ~valid0_o) || (pop3_w && ~valid1_o) || (pop3_w && ~valid2_o) ||
//                        (pop0_w && pop1_w && pop2_w && pop3_w));

integer i;

always @ (posedge clk_i or posedge rst_i)
if (rst_i)
begin
    count_q   <= {(COUNT_W) {1'b0}};
    rd_ptr_q  <= {(ADDR_W) {1'b0}};
    wr_ptr_q  <= {(ADDR_W) {1'b0}};

    for (i = 0; i < DEPTH; i = i + 1) 
    begin
        ram_q[i]         <= {(WIDTH) {1'b0}};
        pc_q[i]          <= 32'b0;
        info0_q[i]       <= {(OPC_INFO_W) {1'b0}};
        info1_q[i]       <= {(OPC_INFO_W) {1'b0}};
        info2_q[i]       <= {(OPC_INFO_W) {1'b0}};
        info3_q[i]       <= {(OPC_INFO_W) {1'b0}};
        valid0_q[i]      <= 1'b0;
        valid1_q[i]      <= 1'b0;
        valid2_q[i]      <= 1'b0;
        valid3_q[i]      <= 1'b0;
    end
end
else if (flush_i)
begin
    count_q   <= {(COUNT_W) {1'b0}};
    rd_ptr_q  <= {(ADDR_W) {1'b0}};
    wr_ptr_q  <= {(ADDR_W) {1'b0}};

    for (i = 0; i < DEPTH; i = i + 1) 
    begin
        info0_q[i]       <= {(OPC_INFO_W) {1'b0}};
        info1_q[i]       <= {(OPC_INFO_W) {1'b0}};
        info2_q[i]       <= {(OPC_INFO_W) {1'b0}};
        info3_q[i]       <= {(OPC_INFO_W) {1'b0}};
        valid0_q[i]      <= 1'b0; // descomentado
        valid1_q[i]      <= 1'b0; // descomentado
        valid2_q[i]      <= 1'b0;
        valid3_q[i]      <= 1'b0;
    end
end
else
begin
    // Push
    if (push_w)
    begin
        ram_q[wr_ptr_q]     <= data_in_i;
        pc_q[wr_ptr_q]      <= pc_in_i;
        info0_q[wr_ptr_q]   <= info0_in_i;
        info1_q[wr_ptr_q]   <= info1_in_i;
        info2_q[wr_ptr_q]   <= info2_in_i;
        info3_q[wr_ptr_q]   <= info3_in_i;
        valid0_q[wr_ptr_q]  <= 1'b1; //sempre valido
        valid1_q[wr_ptr_q]  <= (pred_in_i >= 2'b01); // valido apenas se 2 ou mais instruções
        valid2_q[wr_ptr_q]  <= (pred_in_i >= 2'b10); // valido apenas se 3 ou 4 instruções
        valid3_q[wr_ptr_q]  <= (pred_in_i >= 2'b11); // valido apenas se 4 instruções
        wr_ptr_q            <= wr_ptr_q + 1;
    end

    if (pop0_w)
        valid0_q[rd_ptr_q] <= 1'b0;
    if (pop1_w)
        valid1_q[rd_ptr_q] <= 1'b0;
    if (pop2_w)
        valid2_q[rd_ptr_q] <= 1'b0;
    if (pop3_w)
        valid3_q[rd_ptr_q] <= 1'b0;

    // Both instructions completed
    if (pop_complete_w)
        rd_ptr_q  <= rd_ptr_q + 1;

    if (push_w & ~pop_complete_w)
        count_q <= count_q + 1;
    else if (~push_w & pop_complete_w)
        count_q <= count_q - 1;
end

//-------------------------------------------------------------------
// Combinatorial
//-------------------------------------------------------------------
/* verilator lint_off WIDTH */
assign valid0_o      = (count_q != 0) & valid0_q[rd_ptr_q];
assign valid1_o      = (count_q != 0) & valid1_q[rd_ptr_q];
assign valid2_o      = (count_q != 0) & valid2_q[rd_ptr_q];
assign valid3_o      = (count_q != 0) & valid3_q[rd_ptr_q];
assign accept_o      = (count_q != DEPTH);
/* verilator lint_on WIDTH */

assign pc0_out_o     = {pc_q[rd_ptr_q][31:4],4'b0000};
assign pc1_out_o     = {pc_q[rd_ptr_q][31:4],4'b0100};
assign pc2_out_o     = {pc_q[rd_ptr_q][31:4],4'b1000};
assign pc3_out_o     = {pc_q[rd_ptr_q][31:4],4'b1100};
assign data0_out_o   = ram_q[rd_ptr_q][(WIDTH/4)-1:0];
assign data1_out_o   = ram_q[rd_ptr_q][(WIDTH/2)-1:(WIDTH/4)];
assign data2_out_o   = ram_q[rd_ptr_q][(3*WIDTH/4)-1:(WIDTH/2)];
assign data3_out_o   = ram_q[rd_ptr_q][WIDTH-1:(3*WIDTH/4)];

assign info0_out_o   = info0_q[rd_ptr_q];
assign info1_out_o   = info1_q[rd_ptr_q];
assign info2_out_o   = info2_q[rd_ptr_q];
assign info3_out_o   = info3_q[rd_ptr_q];
endmodule